`timescale 1ns / 100ps

/*

Camera Core (Couple with an architecture-specific wrapper)

Overview

    Camera Core is made of two sub modules and a little glue logic:

    - camera_config    - handles sending the correct I2C commands to get the camera to run
    - i2c_master_core  - handles I2C communication with the camera

    Output is in the form of a pixel stream

    SCL & SDA, being special signals, are finalized in the layers above (architecturally dependent)

    The XCLK (SYSCLK) is special too.  It too is generated by the layers above.

    At this level, the signals should have appropriate names from the datasheet where possible.

Main States

    POWER_OFF

    CONFIGURING - the module is sending all the control signals to the device

    RUNNABLE - the camera is runnable - either running or idle, sending images
        when running, and receptive to commands (like set_origin, etc.)

Configuration

    The camera requires its nReset line to be held low for some number of SYSCLKS.  The FPGA reset
    line is used for this - it is slow to come up after the clock starts.

    As is often the case, finding register values, defaults, etc. is a bit of a Google treasure hunt.

    The registers, default values, etc. are all defined in the camera_config  module.  Those values
    that are configurable by this code (as opposed to being fixed) are presented either as parameters
    or ports.

    After power up, when requested by `configure` the camera is sent the configuration settings.  It then
    waits for the `start` signal to start running.

    While in this configured state, commands like set_window, etc. can be run.

    At this point it sends the RESET and starts running.

Output

    The pixel output from this module is identical to the camera output except a) it is only active
    when the module is running, and b) pclk is replaced by a one clock valid signal.

Hardware

    THe On Semi datasheet is much nicer than the Aptina one.

            |Pin No.|PIN NAME  | TYPE   |DESCRIPTION|
            | - | -            | -      | - |
            | 1 | VCC          | POWER  | 3.3v Power supply |
            | 2 | GND          | Ground | Power ground |
            | 3 | SCL          | Input  | Two-Wire Serial Interface Clock |
            | 4 | SDA(SDATA)   | Bi-directional | Two-Wire Serial Interface Data I/O |
            | 5 | VS(VSYNC)    | Output | Active High: Frame Valid; indicates active frame |
            | 6 | HS(HREF)     | Output | Active High: Line/Data Valid; indicates active pixels |
            | 7 | PCLK         | Output | Pixel Clock output from sensor |
            | 8 | XCLK         | Input  | Master Clock into Sensor (13MHz - 27MHz) |
            | 9 | D9           | Output | Pixel Data Output 9(MSB) |
            | 10| D8           | Output | Pixel Data Output 7(MSB) |
            | 11| D7           | Output | Pixel Data Output 7(MSB) |
            | 12| D6           | Output | Pixel Data Output 6      |
            | 13| D5           | Output | Pixel Data Output 5      |
            | 14| D4           | Output | Pixel Data Output 4      |
            | 15| D3           | Output | Pixel Data Output 3      |
            | 16| D2           | Output | Pixel Data Output 2      |
            | 17| D1           | Output | Pixel Data Output 1      |
            | 18| D0           | Output | Pixel Data Output 0 (LSB)|
            | 19| RST          | Input  | Sensor Reset |
            | 20| PDN(PWDN)    | Input  | |
            | 21| Trigger(EXP) | Input | External trigger output  (confirm Input!?) |
            | 22| LED          | Output | LED Strobe, Exposure indicator |

    - Module requires a SYSCLK (13MHz - 27MHz), halving the 48 seems reasonable.
    - RESET (active low) must be applied for at least 10 SYSCLK cycles after power up
    - STANDBY (active high) must be low
    - Arducam datasheet is wrong about Pins 21 & 22  (they're swapped.  The above is correct)  21 is the trigger.

    Pixel Data

        Simultaneous Master Mode - Continuous frames, exposure happens during the previous frame.  Exposure is indicated
        by LED_Out.  Makes sense.

                        _...__________
            LED_Out   _/              \____________________________________________..._____________________________
                      ___...___        ____________________________________________..._________________________
            Frame              \______/                                                                        \___
                                                  _________         ________                _________
            Line      ___...___|______|__________/         \_______/        \______..._____/         \________|____
                               |      |          |         |       |        |              |         |        |
                       P2      |  V   |    P1    |    A    |   Q   |   A    |   Q       Q  |    A    |   P2   |


                Frame Blanking in this mode may be extended when the exposure time is longer than the frame time

        Snapshot Mode - Exposure is triggered, when complete the frame is sent

                         _
            Exposure  __/ \__..._________________________________________________..._______________________________
                           __...___
            LED_Out   ____/        \_____________________________________________..._______________________________
                                     ____________________________________________...__________________________
            Frame     _______...____/                                                                         \____
                                                _________         ________                _________
            Line      _______...____|__________/         \_______/        \______..._____/         \________|______
                                    |          |         |       |        |              |         |        |
                                    |    P1    |    A    |   Q   |   A    |   Q       Q  |    A    |   P2   |

            V     = Vertical Blanking     = R06
            P1    = Frame Start Blanking  = R05 - 23
            A     = Active Data Time      = R04
            Q     = Horizontal Blanking   = R05
            P2    = Frame End Blanking    = 23 (fixed)

            R     = Rows

            A + Q = Row Time

            F     = Total Frame Time = V + R x ( A + Q )


Issues

    - The busy signal takes a cycle or two to come up (at least 1!), so remember to give it a
      little bit after issuing a command.

    - Probably need a low power mode

    - Is the IDLE vs RUNNING distinction useful?  A way to stop output is probably good, even
      if the camera is still sending

Use



Invocation


Sub Modules

    camera_config
    camera_image

Testing

    Tested in camera_tb.v

    Tested on the Hackaday 2019 Badge (ECP5)

*/

`include "../../pipe/rtl/pipe_defs.v"

module camera_core #(
        parameter Width = 752,
        parameter Height = 482,
        parameter CoordinateWidth = 10,
        parameter BlankingWidth = 16,
        parameter CameraPixelWidth = 10,
        parameter I2CClockCount = 200,
        parameter I2CGapCount = ( 1 << 8 )
    ) (
        input clock,
        input reset,

        // Camera Control
        // input  power_up, // future
        input  configure,
        input  start,
        input  stop,
        // input  power_down, // future

        // Camera Status
        output configuring,
        output error,
        output idle,
        output running,
        output busy,

        // Configuration Commands
        input [CoordinateWidth-1:0] column_start,
        input [CoordinateWidth-1:0] row_start,
        input [CoordinateWidth-1:0] window_width,
        input [CoordinateWidth-1:0] window_height,

        input set_origin,
        input set_window,

        input [BlankingWidth-1:0]   horizontal_blanking,
        input [BlankingWidth-1:0]   vertical_blanking,

        input set_blanking,

        input snapshot_mode,
        input set_snapshot_mode,
        input snapshot,

        // Data Output
        output  out_vs,
        output  out_hs,
        output  out_valid,
        output  [CameraPixelWidth-1:0] out_d,

        // Camera Connections
        output scl_out,
        input  scl_in,
        output sda_out,
        input  sda_in,

        input  vs,
        input  hs,
        input  pclk,

        input  [CameraPixelWidth-1:0] d,

        output rst,
        output pwdn,

        input  led,
        output trigger,

        output [7:0] debug
    );

    // Spec the pipe- a standard 8bit pipe with Start Stop message markers
    localparam I2CPipeSpec = `PS_d8s;
    localparam I2CPipeWidth = `P_w( I2CPipeSpec );
    localparam I2CPipeDataWidth = `P_Data_w( I2CPipeSpec );

    //
    // Control
    //

    reg c_configuring;
    reg c_running;
    reg c_idle;
    reg c_error;

    assign configuring = c_configuring;
    assign running = c_running;
    assign idle = c_idle;

    reg c_rst;
    reg c_pwdn;
    reg c_trigger;

    assign rst = c_rst;
    assign pwdn = c_pwdn;
    assign trigger = c_trigger;

    //
    // I2C Pipe
    //

    wire [I2CPipeWidth-1:0]  config_to_i2c_pipe;
    wire [I2CPipeWidth-1:0]  i2c_to_config_pipe;

    //
    // Camera Config
    //

    reg config_configure;
    reg config_start;
    reg config_stop;
    wire config_running;
    wire config_idle;

    camera_config #(
            .CoordinateWidth( CoordinateWidth ),
            .BlankingWidth( BlankingWidth ),
            .PS( I2CPipeSpec ),
            .I2CGapCount( I2CGapCount )
        ) cam_conf (
            .clock( clock ),
            .reset( reset ),

            .configure( config_configure ),
            .start( config_start ),
            .stop( config_stop ),

            .running( config_running ),
            .idle( config_idle ),
            .busy( busy ),   // direct to the camera_core ports
            .error( error ), // direct to the camera_core ports

            // all window and blanking commands go direct
            .column_start( column_start ),
            .row_start( row_start),
            .window_width( window_width ),
            .window_height( window_height ),

            .set_origin( set_origin ),
            .set_window( set_window ),

            .horizontal_blanking( horizontal_blanking ),
            .vertical_blanking( vertical_blanking ),

            .set_blanking( set_blanking ),

            .snapshot_mode( snapshot_mode ),
            .set_snapshot_mode( set_snapshot_mode ),

            .i2c_pipe_out( config_to_i2c_pipe ),
            .i2c_pipe_in( i2c_to_config_pipe )
        );

    //
    // I2C Master
    //
    // Connected to the Config module via two pipes.
    //
    // Using the Core version here - dragging the architecture-neutral *4* I2C wires all the way out.
    //

    // 8'HB9 is the "READ address"
    // 8'HB8 is the "WRITE address"
    // Actual address without the B0 R/W is 8'H5C
    localparam SlaveAddress = (8'H48);

    i2c_master_core #(
            .PipeSpec( I2CPipeSpec ),
            .ClockCount( I2CClockCount )
        ) i2c_m(
            .clock( clock ),
            .reset( reset ),

            // Set up
            .slave_address( SlaveAddress ),     // slave address is fixed, therefore not sent every time
            .read_count( 9'H1FF ),              // not specified here - in message (-1)
            .operation( 3'H7 ),                 // not specified here - in message (-1)
            .send_address( 1'H0 ),              // no need to pack the address in the return message
            .send_operation( 1'H0 ),            // do return the operation
            .send_write_count( 1'H1 ),          // do return the write count

            .start_operation( 1'H0 ),           // needed only for operations that have no in-pipe config component

            // Pipes in and out
            .pipe_in( config_to_i2c_pipe ),
            .pipe_out( i2c_to_config_pipe ),

            // I2C Lines (in and out broken up to maintain architectural neutrality
            .scl_in( scl_in ),
            .scl_out( scl_out ),
            .sda_out( sda_out ),
            .sda_in( sda_in )

            //.debug( debug )
        );

    //
    // Camera Control
    //

    localparam C_POWERUP = 0,
               C_RESET = 1,
               C_CONFIGURING = 2,
               C_RUNNABLE = 3;

    reg [2:0] c_state;

    always @( posedge clock ) begin

        if ( reset ) begin
            config_start <= 0;
            config_stop <= 0;
            c_running <= 0;
            c_configuring <= 0;
            c_idle <= 0;
            c_rst <= 0;  // device is held in reset
            c_pwdn <= 0;
            c_trigger <= 0;
            c_state <= C_POWERUP;
        end else begin
            case ( c_state )
                C_POWERUP: begin
                        // clear reset
                        c_rst <= 1;
                        c_state <= C_RESET;
                    end
                C_RESET: begin
                        if ( configure ) begin
                            config_configure <= 1;
                            c_configuring <= 1;
                            c_state <= C_CONFIGURING;
                        end
                    end
                C_CONFIGURING: begin
                        config_configure <= 0;
                        if ( error ) begin
                            c_configuring <= 0;
                            c_state <= C_POWERUP;
                        end else begin
                            if ( config_idle ) begin
                                c_configuring <= 0;
                                c_idle <= 1;
                                c_state <= C_RUNNABLE;
                            end
                        end
                    end
                C_RUNNABLE: begin
                        if ( start ) begin
                            c_idle <= 0;
                            c_running <= 1;
                            config_start <= 1;
                            config_stop <= 0;
                        end else begin
                            config_start <= 0;
                            if ( stop ) begin
                                c_idle <= 1;
                                c_running <= 0;
                                config_start <= 0;
                                config_stop <= 1;
                            end else begin
                                config_stop <= 0;
                                if ( snapshot )
                                    c_trigger <= 1;
                                else
                                    c_trigger <= 0;
                            end
                        end
                    end
            endcase
        end

    end

    //
    // Camera Data
    //

    // Ensure two things: data goes out only when the module is in running state, and only full frames go out

    localparam C_OUT_STATE_IDLE = 0,
               C_OUT_STATE_STARTING = 1,
               C_OUT_STATE_RUNNING = 2,
               C_OUT_STATE_STOPPING= 3;

    reg [ 1:0 ] c_out_state;

    reg [ 1:0 ] pclk_history;

    reg [ CameraPixelWidth-1:0 ] c_out_data;

    always @( posedge clock ) begin
        if ( reset ) begin
            c_out_state <= 0;
            c_out_data <= 0;
            pclk_history <= 0;
        end else begin
            pclk_history <= { pclk_history[ 0 ], pclk };
            case ( c_out_state )
                C_OUT_STATE_IDLE:
                    if ( c_running )
                        c_out_state <= C_OUT_STATE_STARTING;
                C_OUT_STATE_STARTING:
                    if ( !vs )
                        c_out_state <= C_OUT_STATE_RUNNING;
                C_OUT_STATE_RUNNING: begin
                        if ( !pclk_history[0] && pclk )
                            c_out_data <= d;
                        if ( !c_running ) begin
                            c_out_state <= C_OUT_STATE_STOPPING;
                        end
                    end
                C_OUT_STATE_STOPPING: begin
                        c_out_data <= 0;
                        if ( !vs )
                            c_out_state <= C_OUT_STATE_IDLE;
                    end
            endcase
        end
    end

    // No output unless c_out_state says so
    wire c_out_running = ( c_out_state == C_OUT_STATE_RUNNING ) || ( c_out_state == C_OUT_STATE_STOPPING );

    assign out_vs    =   ( c_out_running) ?   vs : 0;
    assign out_hs    =   ( c_out_running) ?   hs : 0;
    assign out_valid =   ( c_out_running) ? ( hs && ( pclk_history == 2'B01 ) ) : 0;
    assign out_d     =   ( c_out_running) ?   c_out_data : 0;

endmodule

//
// Camera Config
//
// Takes camera configuration information as parameters, provides initialization sequences
// on its outport designed to connect to the (suitably configured) I2C Master.
//
// Split internally into two levels - the sequencer and the I2C comms io
//
// Address is not sent in the packet, however operation and read size are.  Also write count
// is expected back.
//

module camera_config #(
        parameter CoordinateWidth = 10,
        parameter BlankingWidth = 16,
        parameter PS = `PS_d8s,
        parameter I2CGapCount = (1 << 8)
    ) (
        input clock,
        input reset,

        input  configure,
        input  start,
        input  stop,

        output configuring,
        output running,
        output idle,
        output busy,
        output error,

        input [CoordinateWidth-1:0] column_start,
        input [CoordinateWidth-1:0] row_start,
        input [CoordinateWidth-1:0] window_width,
        input [CoordinateWidth-1:0] window_height,

        input set_origin,
        input set_window,

        input [BlankingWidth-1:0]   horizontal_blanking,
        input [BlankingWidth-1:0]   vertical_blanking,

        input set_blanking,

        input snapshot_mode,
        input set_snapshot_mode,

        inout [`P_w( PS )-1:0] i2c_pipe_in,
        inout [`P_w( PS )-1:0] i2c_pipe_out
    );

    //
    // Camera Registers
    //

    `include "../../drivers/rtl/camera_defs.vh"

    //
    // Output regs
    //

    reg cc_configuring;
    reg cc_idle;
    reg cc_running;
    reg cc_error;
    reg cc_busy;

    reg [CoordinateWidth-1:0] cc_column_start;
    reg [CoordinateWidth-1:0] cc_row_start;
    reg [CoordinateWidth-1:0] cc_window_width;
    reg [CoordinateWidth-1:0] cc_window_height;

    reg [BlankingWidth-1:0]   cc_horizontal_blanking;
    reg [BlankingWidth-1:0]   cc_vertical_blanking;

    reg                       cc_snapshot_mode;

    assign idle = cc_idle;
    assign running = cc_running;
    assign error = cc_error;
    assign busy = cc_busy;

    localparam PipeWidth = `P_w( PS );
    localparam PipeDataWidth = `P_Data_w( PS );

    //
    // Settings
    //

    localparam MaxWidth = 752;
    localparam MaxHeight = 480;
    localparam MinWidth = 48;
    localparam MinHeight = 32;

    localparam ConfigurationResetIndex = 0;
    localparam ConfigurationWindowIndex = 15;
    localparam ConfigurationOriginIndex = 17;
    localparam ConfigurationBlankingIndex = 20;
    localparam ConfigurationSnapshotModeIndex = 23;

    //
    // State Machine
    //

    localparam CC_POWER_OFF     = 0,
               CC_CONNECT       = 1,
               CC_VERSION       = 2,
               CC_CONFIGURE     = 3,
               CC_START         = 4,
               CC_RUNNABLE       = 5;

    reg [2:0]  cc_state;

    // Communication with the I2C SM
    // .. toggle tick to start
    // .. don't mess with the operation details until it's done
    reg        cc_i2c_tick;
    reg        cc_i2c_tock;
    reg        cc_i2c_operation;  // write = 0, read = 1
    reg [7:0]  cc_i2c_register;
    reg [7:0]  cc_i2c_length;
    reg [15:0] cc_i2c_data_in;    // data sent
    reg [15:0] cc_i2c_data_out;   // data returned
    reg [7:0]  cc_i2c_result;     // confirmed length of read or write

    // ...keep these the same as the R/W bit in the I2C standard
    localparam CC_I2C_OPERATION_READ  = 1,
               CC_I2C_OPERATION_WRITE = 0;

    localparam CommsTimerWidth = 26;
    localparam CommsTimerLongCount = I2CGapCount; // During simulation, this needs to be small!  Also not too small.
    localparam CommsTimerShortCount = 10;

    reg [ CommsTimerWidth:0 ] comms_timer;
    wire comms_timer_expired = comms_timer[ CommsTimerWidth ];

    wire       cc_i2c_ready = ( cc_i2c_tick == cc_i2c_tock );
    wire       cc_i2c_busy  = ( cc_i2c_tick != cc_i2c_tock );

    reg [4:0] cc_configuration_index;

    always @( posedge clock ) begin

        if ( reset ) begin
            cc_state <= CC_POWER_OFF;
            cc_i2c_tick <= 0;
            cc_idle <= 0;
            cc_configuring <= 0;
            cc_running <= 0;
            cc_error <= 0;
            cc_busy <= 1;
            cc_i2c_operation <= 0;
            cc_i2c_register <= 0;
            cc_i2c_length <= 0;
            cc_i2c_data_out <= 0;
            cc_configuration_index <= ConfigurationResetIndex;
            comms_timer <= CommsTimerLongCount;
            cc_column_start <= 0;
            cc_row_start <= 0;
            cc_window_width <= 0;
            cc_window_height <= 0;
            cc_horizontal_blanking <= 0;
            cc_vertical_blanking <= 0;
            cc_snapshot_mode <= 0;

        end else begin
            case ( cc_state )
                CC_POWER_OFF: begin // 0
                        // start configuring
                        if ( configure ) begin
                            cc_error <= 0;
                            cc_state <= CC_CONNECT;
                            comms_timer <= CommsTimerLongCount;
                            cc_configuring <= 1;
                            cc_busy <= 1;
                        end
                    end
                CC_CONNECT: begin // 1
                        if ( cc_i2c_ready ) begin
                            if ( comms_timer_expired ) begin
                                cc_i2c_operation <= CC_I2C_OPERATION_READ;
                                cc_i2c_length <= 2;
                                cc_i2c_register <= Register_ChipVersion;
                                cc_i2c_tick <= !cc_i2c_tick;
                                cc_state <= CC_VERSION;
                                comms_timer <= CommsTimerLongCount;
                            end else begin
                                comms_timer <= comms_timer - 1;
                            end
                        end
                    end
                CC_VERSION: begin // 2
                        if ( cc_i2c_ready ) begin
                            if ( comms_timer_expired ) begin
                                if ( ( cc_i2c_result == cc_i2c_length ) && ( ( cc_i2c_data_in == Register_ChipVersion_MT9V022 ) || ( cc_i2c_data_in == Register_ChipVersion_MT9V034 ) ) ) begin
                                    cc_configuration_index <= ConfigurationResetIndex;
                                    cc_state <= CC_CONFIGURE;
                                    cc_i2c_length <= 2;
                                    // comms_timer <= CommsTimerLongCount;
                                end else begin
                                    cc_error <= 1;
                                    cc_state <= CC_POWER_OFF;
                                end
                            end else begin
                                comms_timer <= comms_timer - 1;
                            end
                        end
                    end
                CC_CONFIGURE: begin // 3
                        if ( cc_i2c_ready ) begin
                            if ( comms_timer_expired ) begin
                                if ( ( cc_i2c_result == cc_i2c_length ) ) begin
                                    if ( cc_configuration_register != 0 ) begin
                                        // Do the next register
                                        cc_configuration_index <= cc_configuration_index + 1;
                                        cc_i2c_operation <= CC_I2C_OPERATION_WRITE;
                                        cc_i2c_length <= 2;
                                        cc_i2c_register <= cc_configuration_register;
                                        cc_i2c_data_out <= cc_configuration_data;
                                        cc_i2c_tick <= !cc_i2c_tick;
                                        comms_timer <= CommsTimerLongCount;
                                    end else begin
                                        cc_configuring <= 0;
                                        if ( cc_running || cc_idle ) begin
                                            cc_state <= CC_RUNNABLE;
                                            cc_busy <= 0;
                                        end else begin
                                            cc_i2c_operation <= CC_I2C_OPERATION_WRITE;
                                            cc_i2c_length <= 2;
                                            cc_i2c_register <= Register_Reset;
                                            cc_i2c_data_out <= Register_Reset_LogicReset_Enable;
                                            cc_i2c_tick <= !cc_i2c_tick;
                                            cc_state <= CC_START;
                                        end
                                    end
                                end else begin
                                    cc_error <= 1;
                                    cc_state <= CC_POWER_OFF;
                                end
                            end else begin
                                comms_timer <= comms_timer - 1;
                            end
                        end
                    end
                CC_START: begin // 4
                        if ( cc_i2c_ready ) begin
                            if ( comms_timer_expired ) begin
                                if ( cc_i2c_result == cc_i2c_length ) begin
                                    cc_idle <= 1;
                                    cc_running <= 0;
                                    cc_busy <= 0;
                                    cc_state <= CC_RUNNABLE;
                                end else begin
                                    cc_error <= 1;
                                    cc_state <= CC_POWER_OFF;
                                end
                            end else begin
                                comms_timer <= comms_timer - 1;
                            end
                        end
                    end
                CC_RUNNABLE: begin // 5
                        comms_timer <= CommsTimerLongCount;
                        case ({ start, stop, set_origin, set_window, set_blanking, set_snapshot_mode })
                            { 1'B1, 1'B0, 1'B0, 1'B0, 1'B0, 1'B0}:  begin // start
                                    cc_running <= 1;
                                    cc_idle <= 0;
                                end
                            { 1'B0, 1'B1, 1'B0, 1'B0, 1'B0, 1'B0}:  begin // stop
                                    cc_running <= 0;
                                    cc_idle <= 1;
                                end
                            { 1'B0, 1'B0, 1'B1, 1'B0, 1'B0, 1'B0}:  begin // set_origin
                                    // latch in the values
                                    cc_column_start <= column_start;
                                    cc_row_start <= row_start;
                                    cc_configuration_index <= ConfigurationOriginIndex;
                                    cc_busy <= 1;
                                    cc_state <= CC_CONFIGURE;
                                end
                            { 1'B0, 1'B0, 1'B0, 1'B1, 1'B0, 1'B0}:  begin // set_window
                                    // latch in the values
                                    cc_column_start <= column_start;
                                    cc_row_start <= row_start;
                                    cc_window_height <= window_height;
                                    cc_window_width <= window_width;
                                    cc_configuration_index <= ConfigurationWindowIndex;
                                    cc_busy <= 1;
                                    cc_state <= CC_CONFIGURE;
                                end
                            { 1'B0, 1'B0, 1'B0, 1'B0, 1'B1, 1'B0}:  begin // set_blanking
                                    cc_horizontal_blanking <= horizontal_blanking;
                                    cc_vertical_blanking <= vertical_blanking;
                                    cc_configuration_index <= ConfigurationBlankingIndex;
                                    cc_busy <= 1;
                                    cc_state <= CC_CONFIGURE;
                                end
                            { 1'B0, 1'B0, 1'B0, 1'B0, 1'B0, 1'B1}:  begin // set_snapshot_mode
                                    cc_snapshot_mode <= snapshot_mode;
                                    cc_configuration_index <= ConfigurationSnapshotModeIndex;
                                    cc_busy <= 1;
                                    cc_state <= CC_CONFIGURE;
                                end
                            default:  begin
                                end
                        endcase
                    end
            endcase
        end

    end

    //
    // CONFIGURATION TABLE
    //

    reg [7:0]  cc_configuration_register;
    reg [15:0] cc_configuration_data;

    localparam cc_chip_control_snapshot_mode = ( Register_ChipControl_Default &
                                         ~( Register_ChipControl_SensorOperatingMode_mask << Register_ChipControl_SensorOperatingMode_l ) ) |
                                         ( Register_ChipControl_SensorOperatingMode_Snapshot <<  Register_ChipControl_SensorOperatingMode_l );
    localparam cc_chip_control_master_mode = Register_ChipControl_Default;

    always @(*) begin
        cc_configuration_register = 8'H00;
        cc_configuration_data = 16'H0000;
        case ( cc_configuration_index )
            0: begin cc_configuration_register <= Register_ColumnStart;          cc_configuration_data <= Register_ColumnStart_Default;  end
            1: begin cc_configuration_register <= Register_RowStart;             cc_configuration_data <= Register_RowStart_Default; end
            2: begin cc_configuration_register <= Register_WindowHeight;         cc_configuration_data <= Register_WindowHeight_Default; end
            3: begin cc_configuration_register <= Register_WindowWidth;          cc_configuration_data <= Register_WindowWidth_Default; end
            4: begin cc_configuration_register <= Register_ChipControl;          cc_configuration_data <= Register_ChipControl_Default; end
            5: begin cc_configuration_register <= Register_ReadMode;             cc_configuration_data <= Register_ReadMode_Default_RCFlip; end
            6: begin cc_configuration_register <= Register_HorizontalBlanking;   cc_configuration_data <= Register_HorizontalBlanking_Min; end
            7: begin cc_configuration_register <= Register_VerticalBlanking;     cc_configuration_data <= Register_VerticalBlanking_Min; end
            8: begin cc_configuration_register <= Register_Mystery20;            cc_configuration_data <= Register_Mystery20_NewDefault; end
            9: begin cc_configuration_register <= Register_Mystery24;            cc_configuration_data <= Register_Mystery24_NewDefault; end
           10: begin cc_configuration_register <= Register_Mystery2B;            cc_configuration_data <= Register_Mystery2B_NewDefault; end
           11: begin cc_configuration_register <= Register_Mystery2F;            cc_configuration_data <= Register_Mystery2F_NewDefault; end
           12: begin cc_configuration_register <= 8'H00;                         cc_configuration_data <= 16'H0000; end
           13: begin cc_configuration_register <= 8'H00;                         cc_configuration_data <= 16'H0000; end
           14: begin cc_configuration_register <= 8'H00;                         cc_configuration_data <= 16'H0000; end
           15: begin cc_configuration_register <= Register_WindowHeight;         cc_configuration_data <= cc_window_height; end
           16: begin cc_configuration_register <= Register_WindowWidth;          cc_configuration_data <= cc_window_width; end
           17: begin cc_configuration_register <= Register_ColumnStart;          cc_configuration_data <= cc_column_start; end
           18: begin cc_configuration_register <= Register_RowStart;             cc_configuration_data <= cc_row_start; end
           19: begin cc_configuration_register <= 8'H00;                         cc_configuration_data <= 16'H0000; end
           20: begin cc_configuration_register <= Register_HorizontalBlanking;   cc_configuration_data <= cc_horizontal_blanking; end
           21: begin cc_configuration_register <= Register_VerticalBlanking;     cc_configuration_data <= cc_vertical_blanking; end
           22: begin cc_configuration_register <= 8'H00;                         cc_configuration_data <= 16'H0000; end
           23: begin cc_configuration_register <= Register_ChipControl;          cc_configuration_data <= ( cc_snapshot_mode ) ?  cc_chip_control_snapshot_mode :  cc_chip_control_master_mode; end
           24: begin cc_configuration_register <= 8'H00;                         cc_configuration_data <= 16'H0000; end
        endcase
    end

            // 0: begin cc_configuration_register <= Register_ColumnStart;          cc_configuration_data <= 16'D136;  end
            // 1: begin cc_configuration_register <= Register_RowStart;             cc_configuration_data <= 16'D80; end
            // 2: begin cc_configuration_register <= Register_WindowHeight;         cc_configuration_data <= 16'D320; end
            // 3: begin cc_configuration_register <= Register_WindowWidth;          cc_configuration_data <= 16'D481; end

            //  0: begin cc_configuration_register <= Register_ColumnStart;             cc_configuration_data <= Register_ColumnStart_Default;  end
            //  1 : begin cc_configuration_register <= Register_RowStart;               cc_configuration_data <= Register_RowStart_Default; end
            //  2: begin cc_configuration_register <= Register_WindowHeight;            cc_configuration_data <= Register_WindowHeight_Default; end
            //  3: begin cc_configuration_register <= Register_WindowWidth;             cc_configuration_data <= Register_WindowWidth_Default; end
            //  4: begin cc_configuration_register <= Register_ChipControl;             cc_configuration_data <= Register_ChipControl_Snapshot_Default; end
            //  6: begin cc_configuration_register <= Register_HorizontalBlanking;      cc_configuration_data <= Register_HorizontalBlanking_Min; end
            //  7: begin cc_configuration_register <= Register_VerticalBlanking;        cc_configuration_data <= Register_VerticalBlanking_Min; end
            //  7: begin cc_configuration_register <= Register_VerticalBlanking;        cc_configuration_data <= Register_VerticalBlanking_Default; end
            //  8: begin cc_configuration_register <= 8'H00;                            cc_configuration_data <= 16'H0000; end
            //  9: begin cc_configuration_register <= Register_AecAgcEnable;            cc_configuration_data <= 16'H0000; end
            // 10: begin cc_configuration_register <= Register_CoarseShutterWidthTotal; cc_configuration_data <= 16'H0100; end


    //
    // I2C Comms IO
    //

    // Pipe signals
    reg          i2c_pipe_out_start;
    reg          i2c_pipe_out_stop;
    reg [PipeDataWidth-1:0] i2c_pipe_out_data;
    reg          i2c_pipe_out_valid;
    wire         i2c_pipe_out_ready;

    // Pack (s)tart (s)top (d)ata (v)alid (r)ready into (p)ipe
    p_pack_ssdvrp #( PS ) i2c_out_pack( i2c_pipe_out_start, i2c_pipe_out_stop, i2c_pipe_out_data, i2c_pipe_out_valid, i2c_pipe_out_ready, i2c_pipe_out );

    wire          i2c_pipe_in_start;
    wire          i2c_pipe_in_stop;
    wire [PipeDataWidth-1:0] i2c_pipe_in_data;
    wire          i2c_pipe_in_valid;
    reg           i2c_pipe_in_ready;

    // Unpack (p)ipe into (s)tart (s)top (d)ata (v)alid (r)ready
    p_unpack_pssdvr #( PS ) i2c_in_unpack(  i2c_pipe_in , i2c_pipe_in_start, i2c_pipe_in_stop, i2c_pipe_in_data, i2c_pipe_in_valid, i2c_pipe_in_ready );

    reg [15:0] cc_i2c_data_out_working;

    localparam CC_I2C_IDLE = 0,
               CC_I2C_WRITE_OPERATION = 1,
               CC_I2C_WRITE_REGISTER = 2,
               CC_I2C_WRITE_GET_STATUS = 3,
               CC_I2C_WRITE_DATA = 4,
               CC_I2C_WRITE_DATA_GET_STATUS = 5,
               CC_I2C_READ_OPERATION = 6,
               CC_I2C_READ_SEND_LENGTH = 7,
               CC_I2C_READ_DATA = 8;

    reg [3:0] cc_i2c_state;

    always @( posedge clock ) begin

        if ( reset ) begin
            cc_i2c_state <= CC_I2C_IDLE;
            cc_i2c_tock <= 0;
            i2c_pipe_out_start <= 0;
            i2c_pipe_out_stop <= 0;
            i2c_pipe_out_data <= 0;
            i2c_pipe_out_valid <= 0;
            i2c_pipe_in_ready <= 0;
            cc_i2c_result <= 0;
            cc_i2c_data_in <= 0;
            cc_i2c_data_out_working <= 0;
        end else begin
            case ( cc_i2c_state )
                CC_I2C_IDLE: begin // 0
                        // check for an operation (leave result alone so upper levels can see how it went)
                        if ( cc_i2c_busy ) begin
                            // can start writing the register to the i2c module
                            i2c_pipe_out_start <= 1;
                            i2c_pipe_out_stop <= 0;
                            i2c_pipe_out_data <= CC_I2C_OPERATION_WRITE;
                            i2c_pipe_out_valid <= 1;
                            cc_i2c_state <= CC_I2C_WRITE_OPERATION;
                            cc_i2c_result <= 0;
                            // could test for silly lengths here - they should be 2
                        end
                    end
                CC_I2C_WRITE_OPERATION: begin // 1
                        // was the operation accepted?
                        if ( i2c_pipe_out_ready ) begin
                            i2c_pipe_out_start <= 0;
                            i2c_pipe_out_data <= cc_i2c_register;
                            cc_i2c_state <= CC_I2C_WRITE_REGISTER;
                            // last byte if we're reading or we're writing no bytes
                            i2c_pipe_out_stop <= ( cc_i2c_operation == CC_I2C_OPERATION_READ ) || ( cc_i2c_length == 0 );
                        end
                    end
                CC_I2C_WRITE_REGISTER: begin // 2
                        // was the register accepted?
                        if ( i2c_pipe_out_ready ) begin
                            if ( ( cc_i2c_operation == CC_I2C_OPERATION_READ ) || ( cc_i2c_length == 0 ) ) begin
                                i2c_pipe_out_stop <= 0;
                                i2c_pipe_out_data <= 0;
                                i2c_pipe_out_valid <= 0;
                                i2c_pipe_in_ready <= 1;
                                cc_i2c_state <= CC_I2C_WRITE_GET_STATUS;
                            end else begin
                                // Operation is a non-zero length WRITE
                                // Set up to send the MSB
                                i2c_pipe_out_data <= cc_i2c_data_out[15:8];
                                cc_i2c_data_out_working <= cc_i2c_data_out[ 7:0 ] << 8;
                                cc_i2c_result <= 1;
                                cc_i2c_state <= CC_I2C_WRITE_DATA;
                            end
                        end
                    end
                CC_I2C_WRITE_GET_STATUS: begin // 3
                        if ( i2c_pipe_in_valid && i2c_pipe_in_start ) begin
                            cc_i2c_result <= 0;
                            if ( cc_i2c_operation == CC_I2C_OPERATION_READ ) begin
                                // if reading, we wrote 1 byte (the camera sees 2 bytes, the address and the register)
                                i2c_pipe_in_ready <= 0;
                                if ( i2c_pipe_in_data == 1 ) begin
                                    // now doing the reading operation
                                    i2c_pipe_out_start <= 1;
                                    i2c_pipe_out_stop <= 0;
                                    i2c_pipe_out_data <= CC_I2C_OPERATION_READ;
                                    i2c_pipe_out_valid <= 1;
                                    cc_i2c_state <= CC_I2C_READ_OPERATION;
                                end else begin
                                    cc_i2c_tock = !cc_i2c_tock;
                                    cc_i2c_state <= CC_I2C_IDLE;
                                end
                            end else begin
                                // cc_i2c_state <= CC_I2C_WRITE_DATA;
                                // i2c_pipe_out_data <= cc_i2c_data_out[ 15:8 ];
                                // cc_i2c_data_out_working <= cc_i2c_data_out[ 7:0 ] << 8;
                                // cc_i2c_result <= 1;
                                // i2c_pipe_out_valid <= 1;
                            end
                        end
                    end
                CC_I2C_WRITE_DATA: begin // 4
                        if ( cc_i2c_result < cc_i2c_length ) begin
                            if ( i2c_pipe_out_ready ) begin
                                // next byte
                                i2c_pipe_out_stop <= 1;
                                i2c_pipe_out_data <= cc_i2c_data_out_working[ 15:8 ];
                                cc_i2c_result <= cc_i2c_result + 1;
                            end
                        end else begin
                            if ( i2c_pipe_out_ready ) begin
                                // shut down the out port
                                i2c_pipe_out_data <= 0;
                                i2c_pipe_out_valid <= 0;
                                i2c_pipe_out_stop <= 0;
                                // wait for the report
                                i2c_pipe_in_ready <= 1;
                                cc_i2c_state <= CC_I2C_WRITE_DATA_GET_STATUS;
                            end
                        end
                    end
                CC_I2C_WRITE_DATA_GET_STATUS: begin // 5
                        if ( i2c_pipe_in_valid && i2c_pipe_in_start ) begin
                                cc_i2c_result <= i2c_pipe_in_data - 1;
                                i2c_pipe_in_ready <= 0;
                                cc_i2c_tock = !cc_i2c_tock;
                                cc_i2c_state <= CC_I2C_IDLE;
                        end
                    end

                CC_I2C_READ_OPERATION: begin // 6
                        if ( i2c_pipe_out_ready ) begin
                            // set up to send read length
                            i2c_pipe_out_start <= 0;
                            i2c_pipe_out_data <= 2;
                            i2c_pipe_out_stop <= 1;
                            cc_i2c_result <= 0;
                            cc_i2c_state <= CC_I2C_READ_SEND_LENGTH;
                        end
                    end
                CC_I2C_READ_SEND_LENGTH: begin // 7
                        if ( i2c_pipe_out_ready ) begin
                            // shut the out port down
                            i2c_pipe_out_data <= 0;
                            i2c_pipe_out_valid <= 0;
                            i2c_pipe_out_stop <= 0;
                            // set up to read data
                            cc_i2c_result <= 0;
                            i2c_pipe_in_ready <= 1;
                            cc_i2c_state <= CC_I2C_READ_DATA;
                        end
                    end
                CC_I2C_READ_DATA: begin // 8
                        if ( i2c_pipe_in_valid && ( i2c_pipe_in_start || cc_i2c_result ) ) begin
                            if ( cc_i2c_result == 0 ) begin
                                cc_i2c_data_in[ 15:8 ] = i2c_pipe_in_data;
                                cc_i2c_result <= 1;
                            end else begin
                                cc_i2c_result <= 2;
                                cc_i2c_data_in[ 7:0 ] = i2c_pipe_in_data;
                                i2c_pipe_in_ready <= 0;
                                cc_i2c_tock = !cc_i2c_tock;
                                cc_i2c_state <= CC_I2C_IDLE;
                            end
                        end
                    end
                default: begin
                        // minimal disabling
                        i2c_pipe_in_ready <= 0;
                        i2c_pipe_out_valid <= 0;
                        // should this happen?
                        cc_i2c_tock = !cc_i2c_tock;
                        // back to idle
                        cc_i2c_state <= CC_I2C_IDLE;
                    end
            endcase
        end

    end

endmodule